//Defining the circuit modules
module VerilogTutorials00(
  //Define the I/O ports
  input a,
  output b
);
  //Assigning the wires 
  assign b = a; //Assign output = input
  //The end of this circuit block
endmodule
